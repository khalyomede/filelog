module file_log

pub enum LogSaveMode {
	single
	daily
}
