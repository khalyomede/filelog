// Todo: extract it in its own package

module filelog

pub enum LogSeverity {
	debug
	info
	notice
	warning
	error
	critical
	alert
	emergency
}
