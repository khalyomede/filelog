module filelog

pub enum LogSaveMode {
	single
	daily
}
