// Todo: extract it in its own package

module file_log

pub enum LogSeverity {
	debug
	info
	notice
	warning
	error
	critical
	alert
	emergency
}
